----------------------------------------------------------------------------
-- cmdProc.vhd
----------------------------------------------------------------------------
-- Brief: A command processor skeleton
----------------------------------------------------------------------------
-- Author: Billy Hou
----------------------------------------------------------------------------


library IEEE;
